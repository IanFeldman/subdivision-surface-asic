`timescale 1ns/1ps

module neighbor
(
    input
);

endmodule

