`timescale 1ns/1ps

module tb_subsurf;

endmodule

