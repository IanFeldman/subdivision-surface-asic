`timescale 1ns/1ps

module subsurf;

endmodule

