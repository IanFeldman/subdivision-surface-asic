`timescale 1ns/1ps

module averager;

endmodule

